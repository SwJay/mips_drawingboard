`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:04:14 06/27/2018 
// Design Name: 
// Module Name:    MIO_BUS 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MIO_BUS(input clk,
					input rst,
					input[3:0]BTN,
					input[15:0]SW,
					input mem_w,
					input[31:0]Cpu_data2bus,				//data from CPU
					input[31:0]addr_bus,
					input[31:0]ram_data_out,
					input[15:0]led_out,
					input[31:0]counter_out,
					input counter0_out,
					input counter1_out,
					input counter2_out,
					
					output reg[31:0]Cpu_data4bus,				//write to CPU
					output reg[31:0]ram_data_in,				//from CPU write to Memory
					output reg[11:0]ram_addr,					//Memory Address signals
					output reg data_ram_we,
					output reg GPIOf0000000_we,				//PIOд/SW��
					output reg GPIOe0000000_we,				//�߶�д
					output reg counter_we,						//counterд�ͳ���
					output reg[31:0]Peripheral_in,
					
					output reg vram_we,
					output reg [11:0] vram_data,
					output reg [18:0] vram_addr,
					input [9:0] ps2kb_key
					);	

	reg data_ram_rd, GPIOf0000000_rd, GPIOe0000000_rd, counter_rd, ps2kb_rd;
	wire counter_over; //��������

	always@(posedge clk) begin
		data_ram_we = 0; //����д�ź�
		data_ram_rd = 0; //������ź�
		counter_we = 0; //������д�ź�
		counter_rd = 0; //���������ź�
		GPIOf0000000_we = 0; //�豸1��PIOд�ź�
		GPIOe0000000_we = 0; //��������Counter_xд�ź�
		GPIOf0000000_rd = 0; //�豸3��4��SW�ȶ��ź�
		GPIOe0000000_rd = 0; //�豸2���߶���ʾ��д�ź�
		ram_addr = 10'h0; //�ڴ������ַ��RAM_B��ַ
		ram_data_in = 32'h0; //�ڴ�д���ݣ�RAM_B��������
		Peripheral_in=32'h0; //�������ߣ�CPU���������д������
		ps2kb_rd = 0; //keyborad

		vram_we = 0; //vga
		vram_data = 12'h0;
		vram_addr = 19'h0;
		case(addr_bus[31:28])
		4'h0:begin // data_ram (00000000 - 00000ffc, actually lower 4KB RAM)
				data_ram_we = mem_w;
				ram_addr = addr_bus[13:2];
				ram_data_in = Cpu_data2bus;
				data_ram_rd = ~mem_w;
		end
		4'he:begin // �߶���ʾ�� (e0000000 - efffffff, SSeg7_Dev)
				GPIOe0000000_we = mem_w;
				Peripheral_in = Cpu_data2bus;
				GPIOe0000000_rd = ~mem_w;
		end
		4'hf:begin // PIO (f0000000 - ffffffff0, 8 LEDs & counter, f000004-fffffff4)
				if(addr_bus[2])begin    //counter 
					counter_we = mem_w;
					Peripheral_in = Cpu_data2bus; //write Counter Value 
					counter_rd = ~mem_w;
				end
				else begin     //LED
					GPIOf0000000_we = mem_w;
					Peripheral_in = Cpu_data2bus; //write Counter set & Initialization and light LED
					GPIOf0000000_rd = ~mem_w;
				end
		end
		4'hc:begin // vram
				vram_we = mem_w;
				vram_addr = addr_bus[18:0];
				vram_data = Cpu_data2bus[11:0];
		end
		4'hd:begin // keyborad
				ps2kb_rd = ~mem_w;
		end
		default:begin;end
		
		endcase
	end
	
always @* begin
	Cpu_data4bus = 32'h0;
		casex({data_ram_rd,GPIOe0000000_rd,counter_rd,GPIOf0000000_rd,ps2kb_rd})
			8'b1xxxx:Cpu_data4bus = ram_data_out; //read from RAM
			8'bx1xxx:Cpu_data4bus = counter_out;  //read from Counter
			8'bxx1xx:Cpu_data4bus = counter_out;  //read from Counter
			8'bxxx1x:Cpu_data4bus = {counter0_out,counter1_out,counter2_out,led_out[12:0],SW}; //read from SW & BTN
			8'bxxxx1:Cpu_data4bus = {{22{1'b0}}, ps2kb_key}; //read from keyborad

		endcase
end


endmodule

